module example (x1, x2, x3, x4, z);
    input x1, x2, x3, x4;
    output z;
    wire x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48;
    assign x5 =  x1 &  x1;
    assign x6 =  x5 &  x2;
    assign x7 =  x6 &  x3;
    assign x8 =  x7 &  x4;
    assign x9 =  x1 &  x1;
    assign x10 = ~x9 &  x2;
    assign x11 =  x10 &  x3;
    assign x12 =  x11 &  x4;
    assign x13 = ~x1 & ~x1;
    assign x14 = ~x13 &  x2;
    assign x15 =  x14 &  x3;
    assign x16 =  x15 &  x4;
    assign x17 =  x1 &  x1;
    assign x18 =  x17 &  x2;
    assign x19 = ~x18 &  x3;
    assign x20 =  x19 &  x4;
    assign x21 =  x1 &  x1;
    assign x22 = ~x21 &  x2;
    assign x23 = ~x22 &  x3;
    assign x24 =  x23 &  x4;
    assign x25 = ~x1 & ~x1;
    assign x26 = ~x25 &  x2;
    assign x27 = ~x26 &  x3;
    assign x28 =  x27 &  x4;
    assign x29 =  x1 &  x1;
    assign x30 =  x29 &  x2;
    assign x31 =  x30 &  x3;
    assign x32 = ~x31 &  x4;
    assign x33 = ~x1 & ~x1;
    assign x34 =  x33 &  x2;
    assign x35 = ~x34 &  x3;
    assign x36 = ~x35 &  x4;
    assign x37 =  x1 &  x1;
    assign x38 = ~x37 &  x2;
    assign x39 = ~x38 &  x3;
    assign x40 = ~x39 &  x4;
    assign x41 = ~x8 & ~x12;
    assign x42 =  x41 & ~x16;
    assign x43 =  x42 & ~x20;
    assign x44 =  x43 & ~x24;
    assign x45 =  x44 & ~x28;
    assign x46 =  x45 & ~x32;
    assign x47 =  x46 & ~x36;
    assign x48 =  x47 & ~x40;
    assign z =  x48;
    
endmodule

